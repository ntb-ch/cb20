-- cb20.vhd

-- Generated using ACDS version 13.0sp1 232 at 2020.06.03.16:36:13

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cb20 is
	port (
		clk_clk                                               : in    std_logic                     := '0';             --                                      clk.clk
		reset_reset_n                                         : in    std_logic                     := '0';             --                                    reset.reset_n
		eim_slave_to_avalon_master_0_conduit_end_ioslv_data   : inout std_logic_vector(15 downto 0) := (others => '0'); -- eim_slave_to_avalon_master_0_conduit_end.ioslv_data
		eim_slave_to_avalon_master_0_conduit_end_isl_cs_n     : in    std_logic                     := '0';             --                                         .isl_cs_n
		eim_slave_to_avalon_master_0_conduit_end_isl_oe_n     : in    std_logic                     := '0';             --                                         .isl_oe_n
		eim_slave_to_avalon_master_0_conduit_end_isl_we_n     : in    std_logic                     := '0';             --                                         .isl_we_n
		eim_slave_to_avalon_master_0_conduit_end_osl_data_ack : out   std_logic;                                        --                                         .osl_data_ack
		eim_slave_to_avalon_master_0_conduit_end_islv_address : in    std_logic_vector(15 downto 0) := (others => '0'); --                                         .islv_address
		dacad5668_0_conduit_end_osl_sclk                      : out   std_logic;                                        --                  dacad5668_0_conduit_end.osl_sclk
		dacad5668_0_conduit_end_oslv_Ss                       : out   std_logic;                                        --                                         .oslv_Ss
		dacad5668_0_conduit_end_osl_mosi                      : out   std_logic;                                        --                                         .osl_mosi
		dacad5668_0_conduit_end_osl_LDAC_n                    : out   std_logic;                                        --                                         .osl_LDAC_n
		dacad5668_0_conduit_end_osl_CLR_n                     : out   std_logic;                                        --                                         .osl_CLR_n
		fqd_interface_0_conduit_end_B                         : in    std_logic_vector(7 downto 0)  := (others => '0'); --              fqd_interface_0_conduit_end.B
		fqd_interface_0_conduit_end_A                         : in    std_logic_vector(7 downto 0)  := (others => '0'); --                                         .A
		gpio_block_0_conduit_end_export                       : inout std_logic_vector(8 downto 0)  := (others => '0'); --                 gpio_block_0_conduit_end.export
		pwm_interface_0_conduit_end_export                    : out   std_logic_vector(3 downto 0);                     --              pwm_interface_0_conduit_end.export
		gpio_block_1_conduit_end_export                       : inout std_logic_vector(7 downto 0)  := (others => '0'); --                 gpio_block_1_conduit_end.export
		watchdog_block_0_wd_signals_granted                   : out   std_logic;                                        --              watchdog_block_0_wd_signals.granted
		watchdog_block_0_wd_signals_watchdog_pwm              : out   std_logic;                                        --                                         .watchdog_pwm
		ppwa_block_0_conduit_end_export                       : in    std_logic_vector(1 downto 0)  := (others => '0')  --                 ppwa_block_0_conduit_end.export
	);
end entity cb20;

architecture rtl of cb20 is
	component cb20_altpll_0 is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component cb20_altpll_0;

	component info_device is
		generic (
			unique_id   : std_logic_vector(31 downto 0)  := "00000000000000000000000000000000";
			description : std_logic_vector(223 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
			dev_size    : integer                        := 0
		);
		port (
			isl_clk             : in  std_logic                     := 'X';             -- clk
			isl_reset_n         : in  std_logic                     := 'X';             -- reset_n
			islv_avs_address    : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			isl_avs_read        : in  std_logic                     := 'X';             -- read
			isl_avs_write       : in  std_logic                     := 'X';             -- write
			islv_avs_write_data : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			oslv_avs_read_data  : out std_logic_vector(31 downto 0);                    -- readdata
			osl_avs_waitrequest : out std_logic;                                        -- waitrequest
			islv_avs_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- byteenable
		);
	end component info_device;

	component eim_slave_to_avalon_master is
		generic (
			TRANSFER_WIDTH : integer := 16
		);
		port (
			ioslv_data       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			isl_cs_n         : in    std_logic                     := 'X';             -- export
			isl_oe_n         : in    std_logic                     := 'X';             -- export
			isl_we_n         : in    std_logic                     := 'X';             -- export
			osl_data_ack     : out   std_logic;                                        -- export
			islv_address     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- export
			isl_clk          : in    std_logic                     := 'X';             -- clk
			isl_reset_n      : in    std_logic                     := 'X';             -- reset_n
			islv_readdata    : in    std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			islv_waitrequest : in    std_logic                     := 'X';             -- waitrequest
			oslv_address     : out   std_logic_vector(15 downto 0);                    -- address
			oslv_read        : out   std_logic;                                        -- read
			oslv_write       : out   std_logic;                                        -- write
			oslv_writedata   : out   std_logic_vector(15 downto 0)                     -- writedata
		);
	end component eim_slave_to_avalon_master;

	component avalon_dacad5668_interface is
		generic (
			BASE_CLK           : integer                       := 33000000;
			SCLK_FREQUENCY     : integer                       := 10000000;
			INTERNAL_REFERENCE : std_logic                     := '0';
			UNIQUE_ID          : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			isl_clk             : in  std_logic                     := 'X';             -- clk
			isl_reset_n         : in  std_logic                     := 'X';             -- reset_n
			osl_sclk            : out std_logic;                                        -- export
			oslv_Ss             : out std_logic;                                        -- export
			osl_mosi            : out std_logic;                                        -- export
			osl_LDAC_n          : out std_logic;                                        -- export
			osl_CLR_n           : out std_logic;                                        -- export
			islv_avs_address    : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			isl_avs_read        : in  std_logic                     := 'X';             -- read
			isl_avs_write       : in  std_logic                     := 'X';             -- write
			islv_avs_write_data : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			oslv_avs_read_data  : out std_logic_vector(31 downto 0);                    -- readdata
			osl_avs_waitrequest : out std_logic;                                        -- waitrequest
			islv_avs_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- byteenable
		);
	end component avalon_dacad5668_interface;

	component avalon_fqd_counter_interface is
		generic (
			number_of_fqds : integer                       := 1;
			unique_id      : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			oslv_avs_read_data  : out std_logic_vector(31 downto 0);                    -- readdata
			isl_avs_read        : in  std_logic                     := 'X';             -- read
			isl_avs_write       : in  std_logic                     := 'X';             -- write
			islv_avs_write_data : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			islv_avs_address    : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			osl_avs_waitrequest : out std_logic;                                        -- waitrequest
			islv_avs_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			isl_clk             : in  std_logic                     := 'X';             -- clk
			isl_reset_n         : in  std_logic                     := 'X';             -- reset_n
			islv_enc_B          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			islv_enc_A          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component avalon_fqd_counter_interface;

	component avalon_pwm_interface is
		generic (
			number_of_pwms : integer                       := 1;
			base_clk       : integer                       := 125000000;
			unique_id      : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			oslv_avs_read_data  : out std_logic_vector(31 downto 0);                    -- readdata
			islv_avs_address    : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			isl_avs_read        : in  std_logic                     := 'X';             -- read
			isl_avs_write       : in  std_logic                     := 'X';             -- write
			islv_avs_write_data : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			osl_avs_waitrequest : out std_logic;                                        -- waitrequest
			islv_avs_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			isl_clk             : in  std_logic                     := 'X';             -- clk
			isl_reset_n         : in  std_logic                     := 'X';             -- reset_n
			oslv_pwm            : out std_logic_vector(3 downto 0)                      -- export
		);
	end component avalon_pwm_interface;

	component avalon_watchdog_interface is
		generic (
			base_clk  : integer                       := 125000000;
			unique_id : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			islv_avs_write_data : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			oslv_avs_read_data  : out std_logic_vector(31 downto 0);                    -- readdata
			isl_avs_write       : in  std_logic                     := 'X';             -- write
			isl_avs_read        : in  std_logic                     := 'X';             -- read
			islv_avs_address    : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			osl_avs_waitrequest : out std_logic;                                        -- waitrequest
			islv_avs_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			isl_clk             : in  std_logic                     := 'X';             -- clk
			isl_reset_n         : in  std_logic                     := 'X';             -- reset_n
			osl_granted         : out std_logic;                                        -- export
			osl_watchdog_pwm    : out std_logic                                         -- export
		);
	end component avalon_watchdog_interface;

	component avalon_ppwa_interface is
		generic (
			number_of_ppwas : integer                       := 1;
			base_clk        : integer                       := 125000000;
			unique_id       : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			islv_avs_write_data     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			oslv_avs_read_data      : out std_logic_vector(31 downto 0);                    -- readdata
			islv_avs_address        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			isl_avs_read            : in  std_logic                     := 'X';             -- read
			isl_avs_write           : in  std_logic                     := 'X';             -- write
			osl_avs_waitrequest     : out std_logic;                                        -- waitrequest
			islv_avs_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			isl_clk                 : in  std_logic                     := 'X';             -- clk
			isl_reset_n             : in  std_logic                     := 'X';             -- reset_n
			islv_signals_to_measure : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component avalon_ppwa_interface;

	component altera_merlin_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(16 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(15 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_translator;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(69 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component altera_merlin_slave_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(16 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(87 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(87 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(88 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(88 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_agent;

	component altera_avalon_sc_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(88 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(88 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component altera_avalon_sc_fifo;

	component cb20_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(69 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component cb20_addr_router;

	component cb20_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(87 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(87 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component cb20_id_router;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component cb20_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(69 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(69 downto 0);                    -- data
			src1_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(69 downto 0);                    -- data
			src2_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(69 downto 0);                    -- data
			src3_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(69 downto 0);                    -- data
			src4_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic;                                        -- endofpacket
			src5_ready         : in  std_logic                     := 'X';             -- ready
			src5_valid         : out std_logic;                                        -- valid
			src5_data          : out std_logic_vector(69 downto 0);                    -- data
			src5_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src5_startofpacket : out std_logic;                                        -- startofpacket
			src5_endofpacket   : out std_logic;                                        -- endofpacket
			src6_ready         : in  std_logic                     := 'X';             -- ready
			src6_valid         : out std_logic;                                        -- valid
			src6_data          : out std_logic_vector(69 downto 0);                    -- data
			src6_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src6_startofpacket : out std_logic;                                        -- startofpacket
			src6_endofpacket   : out std_logic;                                        -- endofpacket
			src7_ready         : in  std_logic                     := 'X';             -- ready
			src7_valid         : out std_logic;                                        -- valid
			src7_data          : out std_logic_vector(69 downto 0);                    -- data
			src7_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src7_startofpacket : out std_logic;                                        -- startofpacket
			src7_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component cb20_cmd_xbar_demux;

	component cb20_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(69 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component cb20_rsp_xbar_demux;

	component cb20_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(69 downto 0);                    -- data
			src_channel         : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                        -- ready
			sink5_valid         : in  std_logic                     := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                        -- ready
			sink6_valid         : in  std_logic                     := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready         : out std_logic;                                        -- ready
			sink7_valid         : in  std_logic                     := 'X';             -- valid
			sink7_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink7_data          : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			sink7_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component cb20_rsp_xbar_mux;

	component cb20_info_device_0_avalon_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(4 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cb20_info_device_0_avalon_slave_translator;

	component cb20_gpio_block_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(3 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cb20_gpio_block_0_avalon_slave_0_translator;

	component cb20_pwm_interface_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(5 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component cb20_pwm_interface_0_avalon_slave_0_translator;

	component cb20_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(69 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(87 downto 0);                    -- data
			out_channel          : out std_logic_vector(7 downto 0);                     -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component cb20_width_adapter;

	component cb20_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(87 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(69 downto 0);                    -- data
			out_channel          : out std_logic_vector(7 downto 0);                     -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component cb20_width_adapter_001;

	component cb20_gpio_block_0 is
		generic (
			number_of_gpios : integer                       := 1;
			unique_id       : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			oslv_avs_read_data  : out   std_logic_vector(31 downto 0);                    -- readdata
			islv_avs_address    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			isl_avs_read        : in    std_logic                     := 'X';             -- read
			isl_avs_write       : in    std_logic                     := 'X';             -- write
			osl_avs_waitrequest : out   std_logic;                                        -- waitrequest
			islv_avs_write_data : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			islv_avs_byteenable : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			isl_clk             : in    std_logic                     := 'X';             -- clk
			isl_reset_n         : in    std_logic                     := 'X';             -- reset_n
			oslv_gpios          : inout std_logic_vector(8 downto 0)  := (others => 'X')  -- export
		);
	end component cb20_gpio_block_0;

	component cb20_gpio_block_1 is
		generic (
			number_of_gpios : integer                       := 1;
			unique_id       : std_logic_vector(31 downto 0) := "00000000000000000000000000000000"
		);
		port (
			oslv_avs_read_data  : out   std_logic_vector(31 downto 0);                    -- readdata
			islv_avs_address    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			isl_avs_read        : in    std_logic                     := 'X';             -- read
			isl_avs_write       : in    std_logic                     := 'X';             -- write
			osl_avs_waitrequest : out   std_logic;                                        -- waitrequest
			islv_avs_write_data : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			islv_avs_byteenable : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			isl_clk             : in    std_logic                     := 'X';             -- clk
			isl_reset_n         : in    std_logic                     := 'X';             -- reset_n
			oslv_gpios          : inout std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component cb20_gpio_block_1;

	signal altpll_0_c0_clk                                                                                        : std_logic;                     -- altpll_0:c0 -> [EIM_Slave_to_Avalon_Master_0:isl_clk, EIM_Slave_to_Avalon_Master_0_avalon_master_translator:clk, EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:clk, addr_router:clk, cmd_xbar_demux:clk, dacad5668_0:isl_clk, dacad5668_0_avalon_slave_translator:clk, dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:clk, dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, fqd_interface_0:isl_clk, fqd_interface_0_avalon_slave_0_translator:clk, fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, gpio_block_0:isl_clk, gpio_block_0_avalon_slave_0_translator:clk, gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, gpio_block_1:isl_clk, gpio_block_1_avalon_slave_0_translator:clk, gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, info_device_0:isl_clk, info_device_0_avalon_slave_translator:clk, info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:clk, info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ppwa_block_0:isl_clk, ppwa_block_0_avalon_slave_0_translator:clk, ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pwm_interface_0:isl_clk, pwm_interface_0_avalon_slave_0_translator:clk, pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_mux:clk, rst_controller_001:clk, watchdog_block_0:isl_clk, watchdog_block_0_avalon_slave_0_translator:clk, watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk, width_adapter_010:clk, width_adapter_011:clk, width_adapter_012:clk, width_adapter_013:clk, width_adapter_014:clk, width_adapter_015:clk]
	signal eim_slave_to_avalon_master_0_avalon_master_waitrequest                                                 : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:av_waitrequest -> EIM_Slave_to_Avalon_Master_0:islv_waitrequest
	signal eim_slave_to_avalon_master_0_avalon_master_writedata                                                   : std_logic_vector(15 downto 0); -- EIM_Slave_to_Avalon_Master_0:oslv_writedata -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:av_writedata
	signal eim_slave_to_avalon_master_0_avalon_master_address                                                     : std_logic_vector(15 downto 0); -- EIM_Slave_to_Avalon_Master_0:oslv_address -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:av_address
	signal eim_slave_to_avalon_master_0_avalon_master_write                                                       : std_logic;                     -- EIM_Slave_to_Avalon_Master_0:oslv_write -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:av_write
	signal eim_slave_to_avalon_master_0_avalon_master_read                                                        : std_logic;                     -- EIM_Slave_to_Avalon_Master_0:oslv_read -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:av_read
	signal eim_slave_to_avalon_master_0_avalon_master_readdata                                                    : std_logic_vector(15 downto 0); -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:av_readdata -> EIM_Slave_to_Avalon_Master_0:islv_readdata
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest                                  : std_logic;                     -- info_device_0:osl_avs_waitrequest -> info_device_0_avalon_slave_translator:av_waitrequest
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0); -- info_device_0_avalon_slave_translator:av_writedata -> info_device_0:islv_avs_write_data
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_address                                      : std_logic_vector(4 downto 0);  -- info_device_0_avalon_slave_translator:av_address -> info_device_0:islv_avs_address
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_write                                        : std_logic;                     -- info_device_0_avalon_slave_translator:av_write -> info_device_0:isl_avs_write
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_read                                         : std_logic;                     -- info_device_0_avalon_slave_translator:av_read -> info_device_0:isl_avs_read
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0); -- info_device_0:oslv_avs_read_data -> info_device_0_avalon_slave_translator:av_readdata
	signal info_device_0_avalon_slave_translator_avalon_anti_slave_0_byteenable                                   : std_logic_vector(3 downto 0);  -- info_device_0_avalon_slave_translator:av_byteenable -> info_device_0:islv_avs_byteenable
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest                                    : std_logic;                     -- dacad5668_0:osl_avs_waitrequest -> dacad5668_0_avalon_slave_translator:av_waitrequest
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0); -- dacad5668_0_avalon_slave_translator:av_writedata -> dacad5668_0:islv_avs_write_data
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_address                                        : std_logic_vector(4 downto 0);  -- dacad5668_0_avalon_slave_translator:av_address -> dacad5668_0:islv_avs_address
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_write                                          : std_logic;                     -- dacad5668_0_avalon_slave_translator:av_write -> dacad5668_0:isl_avs_write
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_read                                           : std_logic;                     -- dacad5668_0_avalon_slave_translator:av_read -> dacad5668_0:isl_avs_read
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0); -- dacad5668_0:oslv_avs_read_data -> dacad5668_0_avalon_slave_translator:av_readdata
	signal dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_byteenable                                     : std_logic_vector(3 downto 0);  -- dacad5668_0_avalon_slave_translator:av_byteenable -> dacad5668_0:islv_avs_byteenable
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest                              : std_logic;                     -- fqd_interface_0:osl_avs_waitrequest -> fqd_interface_0_avalon_slave_0_translator:av_waitrequest
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0); -- fqd_interface_0_avalon_slave_0_translator:av_writedata -> fqd_interface_0:islv_avs_write_data
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                  : std_logic_vector(4 downto 0);  -- fqd_interface_0_avalon_slave_0_translator:av_address -> fqd_interface_0:islv_avs_address
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                    : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator:av_write -> fqd_interface_0:isl_avs_write
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                     : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator:av_read -> fqd_interface_0:isl_avs_read
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0); -- fqd_interface_0:oslv_avs_read_data -> fqd_interface_0_avalon_slave_0_translator:av_readdata
	signal fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);  -- fqd_interface_0_avalon_slave_0_translator:av_byteenable -> fqd_interface_0:islv_avs_byteenable
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest                                 : std_logic;                     -- gpio_block_0:osl_avs_waitrequest -> gpio_block_0_avalon_slave_0_translator:av_waitrequest
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0); -- gpio_block_0_avalon_slave_0_translator:av_writedata -> gpio_block_0:islv_avs_write_data
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                     : std_logic_vector(3 downto 0);  -- gpio_block_0_avalon_slave_0_translator:av_address -> gpio_block_0:islv_avs_address
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                       : std_logic;                     -- gpio_block_0_avalon_slave_0_translator:av_write -> gpio_block_0:isl_avs_write
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                        : std_logic;                     -- gpio_block_0_avalon_slave_0_translator:av_read -> gpio_block_0:isl_avs_read
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(31 downto 0); -- gpio_block_0:oslv_avs_read_data -> gpio_block_0_avalon_slave_0_translator:av_readdata
	signal gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                                  : std_logic_vector(3 downto 0);  -- gpio_block_0_avalon_slave_0_translator:av_byteenable -> gpio_block_0:islv_avs_byteenable
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest                              : std_logic;                     -- pwm_interface_0:osl_avs_waitrequest -> pwm_interface_0_avalon_slave_0_translator:av_waitrequest
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0); -- pwm_interface_0_avalon_slave_0_translator:av_writedata -> pwm_interface_0:islv_avs_write_data
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                  : std_logic_vector(5 downto 0);  -- pwm_interface_0_avalon_slave_0_translator:av_address -> pwm_interface_0:islv_avs_address
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                    : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator:av_write -> pwm_interface_0:isl_avs_write
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                     : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator:av_read -> pwm_interface_0:isl_avs_read
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0); -- pwm_interface_0:oslv_avs_read_data -> pwm_interface_0_avalon_slave_0_translator:av_readdata
	signal pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                               : std_logic_vector(3 downto 0);  -- pwm_interface_0_avalon_slave_0_translator:av_byteenable -> pwm_interface_0:islv_avs_byteenable
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest                                 : std_logic;                     -- gpio_block_1:osl_avs_waitrequest -> gpio_block_1_avalon_slave_0_translator:av_waitrequest
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0); -- gpio_block_1_avalon_slave_0_translator:av_writedata -> gpio_block_1:islv_avs_write_data
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_address                                     : std_logic_vector(3 downto 0);  -- gpio_block_1_avalon_slave_0_translator:av_address -> gpio_block_1:islv_avs_address
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_write                                       : std_logic;                     -- gpio_block_1_avalon_slave_0_translator:av_write -> gpio_block_1:isl_avs_write
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_read                                        : std_logic;                     -- gpio_block_1_avalon_slave_0_translator:av_read -> gpio_block_1:isl_avs_read
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(31 downto 0); -- gpio_block_1:oslv_avs_read_data -> gpio_block_1_avalon_slave_0_translator:av_readdata
	signal gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                                  : std_logic_vector(3 downto 0);  -- gpio_block_1_avalon_slave_0_translator:av_byteenable -> gpio_block_1:islv_avs_byteenable
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest                             : std_logic;                     -- watchdog_block_0:osl_avs_waitrequest -> watchdog_block_0_avalon_slave_0_translator:av_waitrequest
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                               : std_logic_vector(31 downto 0); -- watchdog_block_0_avalon_slave_0_translator:av_writedata -> watchdog_block_0:islv_avs_write_data
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                 : std_logic_vector(4 downto 0);  -- watchdog_block_0_avalon_slave_0_translator:av_address -> watchdog_block_0:islv_avs_address
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                   : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator:av_write -> watchdog_block_0:isl_avs_write
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                    : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator:av_read -> watchdog_block_0:isl_avs_read
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                : std_logic_vector(31 downto 0); -- watchdog_block_0:oslv_avs_read_data -> watchdog_block_0_avalon_slave_0_translator:av_readdata
	signal watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                              : std_logic_vector(3 downto 0);  -- watchdog_block_0_avalon_slave_0_translator:av_byteenable -> watchdog_block_0:islv_avs_byteenable
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest                                 : std_logic;                     -- ppwa_block_0:osl_avs_waitrequest -> ppwa_block_0_avalon_slave_0_translator:av_waitrequest
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0); -- ppwa_block_0_avalon_slave_0_translator:av_writedata -> ppwa_block_0:islv_avs_write_data
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                     : std_logic_vector(4 downto 0);  -- ppwa_block_0_avalon_slave_0_translator:av_address -> ppwa_block_0:islv_avs_address
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                       : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator:av_write -> ppwa_block_0:isl_avs_write
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                        : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator:av_read -> ppwa_block_0:isl_avs_read
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(31 downto 0); -- ppwa_block_0:oslv_avs_read_data -> ppwa_block_0_avalon_slave_0_translator:av_readdata
	signal ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                                  : std_logic_vector(3 downto 0);  -- ppwa_block_0_avalon_slave_0_translator:av_byteenable -> ppwa_block_0:islv_avs_byteenable
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_waitrequest            : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_waitrequest
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_burstcount             : std_logic_vector(1 downto 0);  -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_burstcount -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_writedata              : std_logic_vector(15 downto 0); -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_writedata -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_address                : std_logic_vector(16 downto 0); -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_address -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_lock                   : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_lock -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_write                  : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_write -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_read                   : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_read -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdata               : std_logic_vector(15 downto 0); -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_readdata
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_debugaccess            : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_debugaccess -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_byteenable             : std_logic_vector(1 downto 0);  -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_byteenable -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdatavalid          : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator:uav_readdatavalid
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                     -- info_device_0_avalon_slave_translator:uav_waitrequest -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);  -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> info_device_0_avalon_slave_translator:uav_burstcount
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0); -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> info_device_0_avalon_slave_translator:uav_writedata
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(16 downto 0); -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> info_device_0_avalon_slave_translator:uav_address
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> info_device_0_avalon_slave_translator:uav_write
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> info_device_0_avalon_slave_translator:uav_lock
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> info_device_0_avalon_slave_translator:uav_read
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0); -- info_device_0_avalon_slave_translator:uav_readdata -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                     -- info_device_0_avalon_slave_translator:uav_readdatavalid -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> info_device_0_avalon_slave_translator:uav_debugaccess
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);  -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> info_device_0_avalon_slave_translator:uav_byteenable
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(88 downto 0); -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(88 downto 0); -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0); -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                     -- dacad5668_0_avalon_slave_translator:uav_waitrequest -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);  -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dacad5668_0_avalon_slave_translator:uav_burstcount
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0); -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dacad5668_0_avalon_slave_translator:uav_writedata
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(16 downto 0); -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> dacad5668_0_avalon_slave_translator:uav_address
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> dacad5668_0_avalon_slave_translator:uav_write
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dacad5668_0_avalon_slave_translator:uav_lock
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> dacad5668_0_avalon_slave_translator:uav_read
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0); -- dacad5668_0_avalon_slave_translator:uav_readdata -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                     -- dacad5668_0_avalon_slave_translator:uav_readdatavalid -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dacad5668_0_avalon_slave_translator:uav_debugaccess
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);  -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dacad5668_0_avalon_slave_translator:uav_byteenable
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(88 downto 0); -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(88 downto 0); -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0); -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator:uav_waitrequest -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);  -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> fqd_interface_0_avalon_slave_0_translator:uav_burstcount
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0); -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> fqd_interface_0_avalon_slave_0_translator:uav_writedata
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(16 downto 0); -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> fqd_interface_0_avalon_slave_0_translator:uav_address
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> fqd_interface_0_avalon_slave_0_translator:uav_write
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> fqd_interface_0_avalon_slave_0_translator:uav_lock
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> fqd_interface_0_avalon_slave_0_translator:uav_read
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0); -- fqd_interface_0_avalon_slave_0_translator:uav_readdata -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator:uav_readdatavalid -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fqd_interface_0_avalon_slave_0_translator:uav_debugaccess
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);  -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> fqd_interface_0_avalon_slave_0_translator:uav_byteenable
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(88 downto 0); -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(88 downto 0); -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0); -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                     -- gpio_block_0_avalon_slave_0_translator:uav_waitrequest -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);  -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> gpio_block_0_avalon_slave_0_translator:uav_burstcount
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0); -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> gpio_block_0_avalon_slave_0_translator:uav_writedata
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(16 downto 0); -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> gpio_block_0_avalon_slave_0_translator:uav_address
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> gpio_block_0_avalon_slave_0_translator:uav_write
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> gpio_block_0_avalon_slave_0_translator:uav_lock
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> gpio_block_0_avalon_slave_0_translator:uav_read
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0); -- gpio_block_0_avalon_slave_0_translator:uav_readdata -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                     -- gpio_block_0_avalon_slave_0_translator:uav_readdatavalid -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> gpio_block_0_avalon_slave_0_translator:uav_debugaccess
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);  -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> gpio_block_0_avalon_slave_0_translator:uav_byteenable
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(88 downto 0); -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(88 downto 0); -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0); -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator:uav_waitrequest -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);  -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> pwm_interface_0_avalon_slave_0_translator:uav_burstcount
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0); -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> pwm_interface_0_avalon_slave_0_translator:uav_writedata
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(16 downto 0); -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> pwm_interface_0_avalon_slave_0_translator:uav_address
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> pwm_interface_0_avalon_slave_0_translator:uav_write
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> pwm_interface_0_avalon_slave_0_translator:uav_lock
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> pwm_interface_0_avalon_slave_0_translator:uav_read
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0); -- pwm_interface_0_avalon_slave_0_translator:uav_readdata -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator:uav_readdatavalid -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pwm_interface_0_avalon_slave_0_translator:uav_debugaccess
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);  -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> pwm_interface_0_avalon_slave_0_translator:uav_byteenable
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(88 downto 0); -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(88 downto 0); -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0); -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                     -- gpio_block_1_avalon_slave_0_translator:uav_waitrequest -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);  -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> gpio_block_1_avalon_slave_0_translator:uav_burstcount
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0); -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> gpio_block_1_avalon_slave_0_translator:uav_writedata
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(16 downto 0); -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> gpio_block_1_avalon_slave_0_translator:uav_address
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> gpio_block_1_avalon_slave_0_translator:uav_write
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> gpio_block_1_avalon_slave_0_translator:uav_lock
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> gpio_block_1_avalon_slave_0_translator:uav_read
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0); -- gpio_block_1_avalon_slave_0_translator:uav_readdata -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                     -- gpio_block_1_avalon_slave_0_translator:uav_readdatavalid -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> gpio_block_1_avalon_slave_0_translator:uav_debugaccess
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);  -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> gpio_block_1_avalon_slave_0_translator:uav_byteenable
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(88 downto 0); -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(88 downto 0); -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0); -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest               : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator:uav_waitrequest -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                : std_logic_vector(2 downto 0);  -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> watchdog_block_0_avalon_slave_0_translator:uav_burstcount
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                 : std_logic_vector(31 downto 0); -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> watchdog_block_0_avalon_slave_0_translator:uav_writedata
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                   : std_logic_vector(16 downto 0); -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> watchdog_block_0_avalon_slave_0_translator:uav_address
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                     : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> watchdog_block_0_avalon_slave_0_translator:uav_write
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                      : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> watchdog_block_0_avalon_slave_0_translator:uav_lock
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                      : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> watchdog_block_0_avalon_slave_0_translator:uav_read
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                  : std_logic_vector(31 downto 0); -- watchdog_block_0_avalon_slave_0_translator:uav_readdata -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid             : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator:uav_readdatavalid -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess               : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> watchdog_block_0_avalon_slave_0_translator:uav_debugaccess
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                : std_logic_vector(3 downto 0);  -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> watchdog_block_0_avalon_slave_0_translator:uav_byteenable
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket        : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid              : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket      : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data               : std_logic_vector(88 downto 0); -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready              : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket     : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid           : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket   : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data            : std_logic_vector(88 downto 0); -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready           : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid         : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data          : std_logic_vector(33 downto 0); -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready         : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator:uav_waitrequest -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);  -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> ppwa_block_0_avalon_slave_0_translator:uav_burstcount
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0); -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> ppwa_block_0_avalon_slave_0_translator:uav_writedata
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(16 downto 0); -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> ppwa_block_0_avalon_slave_0_translator:uav_address
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> ppwa_block_0_avalon_slave_0_translator:uav_write
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> ppwa_block_0_avalon_slave_0_translator:uav_lock
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> ppwa_block_0_avalon_slave_0_translator:uav_read
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0); -- ppwa_block_0_avalon_slave_0_translator:uav_readdata -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator:uav_readdatavalid -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ppwa_block_0_avalon_slave_0_translator:uav_debugaccess
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);  -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> ppwa_block_0_avalon_slave_0_translator:uav_byteenable
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(88 downto 0); -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(88 downto 0); -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0); -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket   : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid         : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data          : std_logic_vector(69 downto 0); -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready         : std_logic;                     -- addr_router:sink_ready -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(87 downto 0); -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                     -- id_router:sink_ready -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(87 downto 0); -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                     -- id_router_001:sink_ready -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(87 downto 0); -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                     -- id_router_002:sink_ready -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(87 downto 0); -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                     -- id_router_003:sink_ready -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(87 downto 0); -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                     -- id_router_004:sink_ready -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(87 downto 0); -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                     -- id_router_005:sink_ready -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket               : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                     : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket             : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                      : std_logic_vector(87 downto 0); -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                     : std_logic;                     -- id_router_006:sink_ready -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(87 downto 0); -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                     -- id_router_007:sink_ready -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal rst_controller_reset_out_reset                                                                         : std_logic;                     -- rst_controller:reset_out -> altpll_0:reset
	signal rst_controller_001_reset_out_reset                                                                     : std_logic;                     -- rst_controller_001:reset_out -> [EIM_Slave_to_Avalon_Master_0_avalon_master_translator:reset, EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:reset, addr_router:reset, cmd_xbar_demux:reset, dacad5668_0_avalon_slave_translator:reset, dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fqd_interface_0_avalon_slave_0_translator:reset, fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, gpio_block_0_avalon_slave_0_translator:reset, gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, gpio_block_1_avalon_slave_0_translator:reset, gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, info_device_0_avalon_slave_translator:reset, info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ppwa_block_0_avalon_slave_0_translator:reset, ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pwm_interface_0_avalon_slave_0_translator:reset, pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_mux:reset, rst_controller_001_reset_out_reset:in, watchdog_block_0_avalon_slave_0_translator:reset, watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset, width_adapter_012:reset, width_adapter_013:reset, width_adapter_014:reset, width_adapter_015:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src0_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_src0_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src0_data -> width_adapter:in_data
	signal cmd_xbar_demux_src0_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src0_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_src1_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src1_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src1_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src1_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_src1_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src1_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_src1_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src1_channel -> width_adapter_002:in_channel
	signal cmd_xbar_demux_src2_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src2_endofpacket -> width_adapter_004:in_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src2_valid -> width_adapter_004:in_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src2_startofpacket -> width_adapter_004:in_startofpacket
	signal cmd_xbar_demux_src2_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src2_data -> width_adapter_004:in_data
	signal cmd_xbar_demux_src2_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src2_channel -> width_adapter_004:in_channel
	signal cmd_xbar_demux_src3_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src3_endofpacket -> width_adapter_006:in_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src3_valid -> width_adapter_006:in_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src3_startofpacket -> width_adapter_006:in_startofpacket
	signal cmd_xbar_demux_src3_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src3_data -> width_adapter_006:in_data
	signal cmd_xbar_demux_src3_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src3_channel -> width_adapter_006:in_channel
	signal cmd_xbar_demux_src4_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src4_endofpacket -> width_adapter_008:in_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src4_valid -> width_adapter_008:in_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src4_startofpacket -> width_adapter_008:in_startofpacket
	signal cmd_xbar_demux_src4_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src4_data -> width_adapter_008:in_data
	signal cmd_xbar_demux_src4_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src4_channel -> width_adapter_008:in_channel
	signal cmd_xbar_demux_src5_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src5_endofpacket -> width_adapter_010:in_endofpacket
	signal cmd_xbar_demux_src5_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src5_valid -> width_adapter_010:in_valid
	signal cmd_xbar_demux_src5_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src5_startofpacket -> width_adapter_010:in_startofpacket
	signal cmd_xbar_demux_src5_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src5_data -> width_adapter_010:in_data
	signal cmd_xbar_demux_src5_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src5_channel -> width_adapter_010:in_channel
	signal cmd_xbar_demux_src6_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src6_endofpacket -> width_adapter_012:in_endofpacket
	signal cmd_xbar_demux_src6_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src6_valid -> width_adapter_012:in_valid
	signal cmd_xbar_demux_src6_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src6_startofpacket -> width_adapter_012:in_startofpacket
	signal cmd_xbar_demux_src6_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src6_data -> width_adapter_012:in_data
	signal cmd_xbar_demux_src6_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src6_channel -> width_adapter_012:in_channel
	signal cmd_xbar_demux_src7_endofpacket                                                                        : std_logic;                     -- cmd_xbar_demux:src7_endofpacket -> width_adapter_014:in_endofpacket
	signal cmd_xbar_demux_src7_valid                                                                              : std_logic;                     -- cmd_xbar_demux:src7_valid -> width_adapter_014:in_valid
	signal cmd_xbar_demux_src7_startofpacket                                                                      : std_logic;                     -- cmd_xbar_demux:src7_startofpacket -> width_adapter_014:in_startofpacket
	signal cmd_xbar_demux_src7_data                                                                               : std_logic_vector(69 downto 0); -- cmd_xbar_demux:src7_data -> width_adapter_014:in_data
	signal cmd_xbar_demux_src7_channel                                                                            : std_logic_vector(7 downto 0);  -- cmd_xbar_demux:src7_channel -> width_adapter_014:in_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                        : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                              : std_logic;                     -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                      : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                               : std_logic_vector(69 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                            : std_logic_vector(7 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                              : std_logic;                     -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                    : std_logic;                     -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                          : std_logic;                     -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                  : std_logic;                     -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                           : std_logic_vector(69 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                        : std_logic_vector(7 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                          : std_logic;                     -- rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal addr_router_src_endofpacket                                                                            : std_logic;                     -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                  : std_logic;                     -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                          : std_logic;                     -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                   : std_logic_vector(69 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                : std_logic_vector(7 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                  : std_logic;                     -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                           : std_logic;                     -- rsp_xbar_mux:src_endofpacket -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                 : std_logic;                     -- rsp_xbar_mux:src_valid -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                         : std_logic;                     -- rsp_xbar_mux:src_startofpacket -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                  : std_logic_vector(69 downto 0); -- rsp_xbar_mux:src_data -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                               : std_logic_vector(7 downto 0);  -- rsp_xbar_mux:src_channel -> EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                 : std_logic;                     -- EIM_Slave_to_Avalon_Master_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal cmd_xbar_demux_src0_ready                                                                              : std_logic;                     -- width_adapter:in_ready -> cmd_xbar_demux:src0_ready
	signal width_adapter_src_endofpacket                                                                          : std_logic;                     -- width_adapter:out_endofpacket -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_src_valid                                                                                : std_logic;                     -- width_adapter:out_valid -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_src_startofpacket                                                                        : std_logic;                     -- width_adapter:out_startofpacket -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_src_data                                                                                 : std_logic_vector(87 downto 0); -- width_adapter:out_data -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_src_ready                                                                                : std_logic;                     -- info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                              : std_logic_vector(7 downto 0);  -- width_adapter:out_channel -> info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_src_endofpacket                                                                              : std_logic;                     -- id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_src_valid                                                                                    : std_logic;                     -- id_router:src_valid -> width_adapter_001:in_valid
	signal id_router_src_startofpacket                                                                            : std_logic;                     -- id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_src_data                                                                                     : std_logic_vector(87 downto 0); -- id_router:src_data -> width_adapter_001:in_data
	signal id_router_src_channel                                                                                  : std_logic_vector(7 downto 0);  -- id_router:src_channel -> width_adapter_001:in_channel
	signal id_router_src_ready                                                                                    : std_logic;                     -- width_adapter_001:in_ready -> id_router:src_ready
	signal width_adapter_001_src_endofpacket                                                                      : std_logic;                     -- width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal width_adapter_001_src_valid                                                                            : std_logic;                     -- width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	signal width_adapter_001_src_startofpacket                                                                    : std_logic;                     -- width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal width_adapter_001_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	signal width_adapter_001_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel
	signal cmd_xbar_demux_src1_ready                                                                              : std_logic;                     -- width_adapter_002:in_ready -> cmd_xbar_demux:src1_ready
	signal width_adapter_002_src_endofpacket                                                                      : std_logic;                     -- width_adapter_002:out_endofpacket -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_002_src_valid                                                                            : std_logic;                     -- width_adapter_002:out_valid -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_002_src_startofpacket                                                                    : std_logic;                     -- width_adapter_002:out_startofpacket -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_002_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_002:out_data -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_002_src_ready                                                                            : std_logic;                     -- dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_002:out_channel -> dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_001_src_endofpacket                                                                          : std_logic;                     -- id_router_001:src_endofpacket -> width_adapter_003:in_endofpacket
	signal id_router_001_src_valid                                                                                : std_logic;                     -- id_router_001:src_valid -> width_adapter_003:in_valid
	signal id_router_001_src_startofpacket                                                                        : std_logic;                     -- id_router_001:src_startofpacket -> width_adapter_003:in_startofpacket
	signal id_router_001_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_001:src_data -> width_adapter_003:in_data
	signal id_router_001_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_001:src_channel -> width_adapter_003:in_channel
	signal id_router_001_src_ready                                                                                : std_logic;                     -- width_adapter_003:in_ready -> id_router_001:src_ready
	signal width_adapter_003_src_endofpacket                                                                      : std_logic;                     -- width_adapter_003:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal width_adapter_003_src_valid                                                                            : std_logic;                     -- width_adapter_003:out_valid -> rsp_xbar_demux_001:sink_valid
	signal width_adapter_003_src_startofpacket                                                                    : std_logic;                     -- width_adapter_003:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal width_adapter_003_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_003:out_data -> rsp_xbar_demux_001:sink_data
	signal width_adapter_003_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_001:sink_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_003:out_channel -> rsp_xbar_demux_001:sink_channel
	signal cmd_xbar_demux_src2_ready                                                                              : std_logic;                     -- width_adapter_004:in_ready -> cmd_xbar_demux:src2_ready
	signal width_adapter_004_src_endofpacket                                                                      : std_logic;                     -- width_adapter_004:out_endofpacket -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_004_src_valid                                                                            : std_logic;                     -- width_adapter_004:out_valid -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_004_src_startofpacket                                                                    : std_logic;                     -- width_adapter_004:out_startofpacket -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_004_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_004:out_data -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_004_src_ready                                                                            : std_logic;                     -- fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_004:out_ready
	signal width_adapter_004_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_004:out_channel -> fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_002_src_endofpacket                                                                          : std_logic;                     -- id_router_002:src_endofpacket -> width_adapter_005:in_endofpacket
	signal id_router_002_src_valid                                                                                : std_logic;                     -- id_router_002:src_valid -> width_adapter_005:in_valid
	signal id_router_002_src_startofpacket                                                                        : std_logic;                     -- id_router_002:src_startofpacket -> width_adapter_005:in_startofpacket
	signal id_router_002_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_002:src_data -> width_adapter_005:in_data
	signal id_router_002_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_002:src_channel -> width_adapter_005:in_channel
	signal id_router_002_src_ready                                                                                : std_logic;                     -- width_adapter_005:in_ready -> id_router_002:src_ready
	signal width_adapter_005_src_endofpacket                                                                      : std_logic;                     -- width_adapter_005:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal width_adapter_005_src_valid                                                                            : std_logic;                     -- width_adapter_005:out_valid -> rsp_xbar_demux_002:sink_valid
	signal width_adapter_005_src_startofpacket                                                                    : std_logic;                     -- width_adapter_005:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal width_adapter_005_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_005:out_data -> rsp_xbar_demux_002:sink_data
	signal width_adapter_005_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_002:sink_ready -> width_adapter_005:out_ready
	signal width_adapter_005_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_005:out_channel -> rsp_xbar_demux_002:sink_channel
	signal cmd_xbar_demux_src3_ready                                                                              : std_logic;                     -- width_adapter_006:in_ready -> cmd_xbar_demux:src3_ready
	signal width_adapter_006_src_endofpacket                                                                      : std_logic;                     -- width_adapter_006:out_endofpacket -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_006_src_valid                                                                            : std_logic;                     -- width_adapter_006:out_valid -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_006_src_startofpacket                                                                    : std_logic;                     -- width_adapter_006:out_startofpacket -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_006_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_006:out_data -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_006_src_ready                                                                            : std_logic;                     -- gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_006:out_ready
	signal width_adapter_006_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_006:out_channel -> gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_003_src_endofpacket                                                                          : std_logic;                     -- id_router_003:src_endofpacket -> width_adapter_007:in_endofpacket
	signal id_router_003_src_valid                                                                                : std_logic;                     -- id_router_003:src_valid -> width_adapter_007:in_valid
	signal id_router_003_src_startofpacket                                                                        : std_logic;                     -- id_router_003:src_startofpacket -> width_adapter_007:in_startofpacket
	signal id_router_003_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_003:src_data -> width_adapter_007:in_data
	signal id_router_003_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_003:src_channel -> width_adapter_007:in_channel
	signal id_router_003_src_ready                                                                                : std_logic;                     -- width_adapter_007:in_ready -> id_router_003:src_ready
	signal width_adapter_007_src_endofpacket                                                                      : std_logic;                     -- width_adapter_007:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal width_adapter_007_src_valid                                                                            : std_logic;                     -- width_adapter_007:out_valid -> rsp_xbar_demux_003:sink_valid
	signal width_adapter_007_src_startofpacket                                                                    : std_logic;                     -- width_adapter_007:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal width_adapter_007_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_007:out_data -> rsp_xbar_demux_003:sink_data
	signal width_adapter_007_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_003:sink_ready -> width_adapter_007:out_ready
	signal width_adapter_007_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_007:out_channel -> rsp_xbar_demux_003:sink_channel
	signal cmd_xbar_demux_src4_ready                                                                              : std_logic;                     -- width_adapter_008:in_ready -> cmd_xbar_demux:src4_ready
	signal width_adapter_008_src_endofpacket                                                                      : std_logic;                     -- width_adapter_008:out_endofpacket -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_008_src_valid                                                                            : std_logic;                     -- width_adapter_008:out_valid -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_008_src_startofpacket                                                                    : std_logic;                     -- width_adapter_008:out_startofpacket -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_008_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_008:out_data -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_008_src_ready                                                                            : std_logic;                     -- pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_008:out_ready
	signal width_adapter_008_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_008:out_channel -> pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_004_src_endofpacket                                                                          : std_logic;                     -- id_router_004:src_endofpacket -> width_adapter_009:in_endofpacket
	signal id_router_004_src_valid                                                                                : std_logic;                     -- id_router_004:src_valid -> width_adapter_009:in_valid
	signal id_router_004_src_startofpacket                                                                        : std_logic;                     -- id_router_004:src_startofpacket -> width_adapter_009:in_startofpacket
	signal id_router_004_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_004:src_data -> width_adapter_009:in_data
	signal id_router_004_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_004:src_channel -> width_adapter_009:in_channel
	signal id_router_004_src_ready                                                                                : std_logic;                     -- width_adapter_009:in_ready -> id_router_004:src_ready
	signal width_adapter_009_src_endofpacket                                                                      : std_logic;                     -- width_adapter_009:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal width_adapter_009_src_valid                                                                            : std_logic;                     -- width_adapter_009:out_valid -> rsp_xbar_demux_004:sink_valid
	signal width_adapter_009_src_startofpacket                                                                    : std_logic;                     -- width_adapter_009:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal width_adapter_009_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_009:out_data -> rsp_xbar_demux_004:sink_data
	signal width_adapter_009_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_004:sink_ready -> width_adapter_009:out_ready
	signal width_adapter_009_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_009:out_channel -> rsp_xbar_demux_004:sink_channel
	signal cmd_xbar_demux_src5_ready                                                                              : std_logic;                     -- width_adapter_010:in_ready -> cmd_xbar_demux:src5_ready
	signal width_adapter_010_src_endofpacket                                                                      : std_logic;                     -- width_adapter_010:out_endofpacket -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_010_src_valid                                                                            : std_logic;                     -- width_adapter_010:out_valid -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_010_src_startofpacket                                                                    : std_logic;                     -- width_adapter_010:out_startofpacket -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_010_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_010:out_data -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_010_src_ready                                                                            : std_logic;                     -- gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_010:out_ready
	signal width_adapter_010_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_010:out_channel -> gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_005_src_endofpacket                                                                          : std_logic;                     -- id_router_005:src_endofpacket -> width_adapter_011:in_endofpacket
	signal id_router_005_src_valid                                                                                : std_logic;                     -- id_router_005:src_valid -> width_adapter_011:in_valid
	signal id_router_005_src_startofpacket                                                                        : std_logic;                     -- id_router_005:src_startofpacket -> width_adapter_011:in_startofpacket
	signal id_router_005_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_005:src_data -> width_adapter_011:in_data
	signal id_router_005_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_005:src_channel -> width_adapter_011:in_channel
	signal id_router_005_src_ready                                                                                : std_logic;                     -- width_adapter_011:in_ready -> id_router_005:src_ready
	signal width_adapter_011_src_endofpacket                                                                      : std_logic;                     -- width_adapter_011:out_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal width_adapter_011_src_valid                                                                            : std_logic;                     -- width_adapter_011:out_valid -> rsp_xbar_demux_005:sink_valid
	signal width_adapter_011_src_startofpacket                                                                    : std_logic;                     -- width_adapter_011:out_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal width_adapter_011_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_011:out_data -> rsp_xbar_demux_005:sink_data
	signal width_adapter_011_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_005:sink_ready -> width_adapter_011:out_ready
	signal width_adapter_011_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_011:out_channel -> rsp_xbar_demux_005:sink_channel
	signal cmd_xbar_demux_src6_ready                                                                              : std_logic;                     -- width_adapter_012:in_ready -> cmd_xbar_demux:src6_ready
	signal width_adapter_012_src_endofpacket                                                                      : std_logic;                     -- width_adapter_012:out_endofpacket -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_012_src_valid                                                                            : std_logic;                     -- width_adapter_012:out_valid -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_012_src_startofpacket                                                                    : std_logic;                     -- width_adapter_012:out_startofpacket -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_012_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_012:out_data -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_012_src_ready                                                                            : std_logic;                     -- watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_012:out_ready
	signal width_adapter_012_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_012:out_channel -> watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_006_src_endofpacket                                                                          : std_logic;                     -- id_router_006:src_endofpacket -> width_adapter_013:in_endofpacket
	signal id_router_006_src_valid                                                                                : std_logic;                     -- id_router_006:src_valid -> width_adapter_013:in_valid
	signal id_router_006_src_startofpacket                                                                        : std_logic;                     -- id_router_006:src_startofpacket -> width_adapter_013:in_startofpacket
	signal id_router_006_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_006:src_data -> width_adapter_013:in_data
	signal id_router_006_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_006:src_channel -> width_adapter_013:in_channel
	signal id_router_006_src_ready                                                                                : std_logic;                     -- width_adapter_013:in_ready -> id_router_006:src_ready
	signal width_adapter_013_src_endofpacket                                                                      : std_logic;                     -- width_adapter_013:out_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal width_adapter_013_src_valid                                                                            : std_logic;                     -- width_adapter_013:out_valid -> rsp_xbar_demux_006:sink_valid
	signal width_adapter_013_src_startofpacket                                                                    : std_logic;                     -- width_adapter_013:out_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal width_adapter_013_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_013:out_data -> rsp_xbar_demux_006:sink_data
	signal width_adapter_013_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_006:sink_ready -> width_adapter_013:out_ready
	signal width_adapter_013_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_013:out_channel -> rsp_xbar_demux_006:sink_channel
	signal cmd_xbar_demux_src7_ready                                                                              : std_logic;                     -- width_adapter_014:in_ready -> cmd_xbar_demux:src7_ready
	signal width_adapter_014_src_endofpacket                                                                      : std_logic;                     -- width_adapter_014:out_endofpacket -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_014_src_valid                                                                            : std_logic;                     -- width_adapter_014:out_valid -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_014_src_startofpacket                                                                    : std_logic;                     -- width_adapter_014:out_startofpacket -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_014_src_data                                                                             : std_logic_vector(87 downto 0); -- width_adapter_014:out_data -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_014_src_ready                                                                            : std_logic;                     -- ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_014:out_ready
	signal width_adapter_014_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_014:out_channel -> ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_007_src_endofpacket                                                                          : std_logic;                     -- id_router_007:src_endofpacket -> width_adapter_015:in_endofpacket
	signal id_router_007_src_valid                                                                                : std_logic;                     -- id_router_007:src_valid -> width_adapter_015:in_valid
	signal id_router_007_src_startofpacket                                                                        : std_logic;                     -- id_router_007:src_startofpacket -> width_adapter_015:in_startofpacket
	signal id_router_007_src_data                                                                                 : std_logic_vector(87 downto 0); -- id_router_007:src_data -> width_adapter_015:in_data
	signal id_router_007_src_channel                                                                              : std_logic_vector(7 downto 0);  -- id_router_007:src_channel -> width_adapter_015:in_channel
	signal id_router_007_src_ready                                                                                : std_logic;                     -- width_adapter_015:in_ready -> id_router_007:src_ready
	signal width_adapter_015_src_endofpacket                                                                      : std_logic;                     -- width_adapter_015:out_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal width_adapter_015_src_valid                                                                            : std_logic;                     -- width_adapter_015:out_valid -> rsp_xbar_demux_007:sink_valid
	signal width_adapter_015_src_startofpacket                                                                    : std_logic;                     -- width_adapter_015:out_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal width_adapter_015_src_data                                                                             : std_logic_vector(69 downto 0); -- width_adapter_015:out_data -> rsp_xbar_demux_007:sink_data
	signal width_adapter_015_src_ready                                                                            : std_logic;                     -- rsp_xbar_demux_007:sink_ready -> width_adapter_015:out_ready
	signal width_adapter_015_src_channel                                                                          : std_logic_vector(7 downto 0);  -- width_adapter_015:out_channel -> rsp_xbar_demux_007:sink_channel
	signal reset_reset_n_ports_inv                                                                                : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                                                           : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [EIM_Slave_to_Avalon_Master_0:isl_reset_n, dacad5668_0:isl_reset_n, fqd_interface_0:isl_reset_n, gpio_block_0:isl_reset_n, gpio_block_1:isl_reset_n, info_device_0:isl_reset_n, ppwa_block_0:isl_reset_n, pwm_interface_0:isl_reset_n, watchdog_block_0:isl_reset_n]

begin

	altpll_0 : component cb20_altpll_0
		port map (
			clk       => clk_clk,                        --       inclk_interface.clk
			reset     => rst_controller_reset_out_reset, -- inclk_interface_reset.reset
			read      => open,                           --             pll_slave.read
			write     => open,                           --                      .write
			address   => open,                           --                      .address
			readdata  => open,                           --                      .readdata
			writedata => open,                           --                      .writedata
			c0        => altpll_0_c0_clk,                --                    c0.clk
			areset    => open,                           --        areset_conduit.export
			locked    => open,                           --        locked_conduit.export
			phasedone => open                            --     phasedone_conduit.export
		);

	info_device_0 : component info_device
		generic map (
			unique_id   => "00010010011100000000000000000001",
			description => "01100011011000100011001000110000001000000111011101101001011101000110100000100000011101110110010001110100001011000010000000110010001110000010111000110101001011100011001000110000001100100011000000000000000000000000000000000000",
			dev_size    => 1024
		)
		port map (
			isl_clk             => altpll_0_c0_clk,                                                       --   clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                          --   reset_sink.reset_n
			islv_avs_address    => info_device_0_avalon_slave_translator_avalon_anti_slave_0_address,     -- avalon_slave.address
			isl_avs_read        => info_device_0_avalon_slave_translator_avalon_anti_slave_0_read,        --             .read
			isl_avs_write       => info_device_0_avalon_slave_translator_avalon_anti_slave_0_write,       --             .write
			islv_avs_write_data => info_device_0_avalon_slave_translator_avalon_anti_slave_0_writedata,   --             .writedata
			oslv_avs_read_data  => info_device_0_avalon_slave_translator_avalon_anti_slave_0_readdata,    --             .readdata
			osl_avs_waitrequest => info_device_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest, --             .waitrequest
			islv_avs_byteenable => info_device_0_avalon_slave_translator_avalon_anti_slave_0_byteenable   --             .byteenable
		);

	eim_slave_to_avalon_master_0 : component eim_slave_to_avalon_master
		generic map (
			TRANSFER_WIDTH => 16
		)
		port map (
			ioslv_data       => eim_slave_to_avalon_master_0_conduit_end_ioslv_data,    --   conduit_end.export
			isl_cs_n         => eim_slave_to_avalon_master_0_conduit_end_isl_cs_n,      --              .export
			isl_oe_n         => eim_slave_to_avalon_master_0_conduit_end_isl_oe_n,      --              .export
			isl_we_n         => eim_slave_to_avalon_master_0_conduit_end_isl_we_n,      --              .export
			osl_data_ack     => eim_slave_to_avalon_master_0_conduit_end_osl_data_ack,  --              .export
			islv_address     => eim_slave_to_avalon_master_0_conduit_end_islv_address,  --              .export
			isl_clk          => altpll_0_c0_clk,                                        --    clock_sink.clk
			isl_reset_n      => rst_controller_001_reset_out_reset_ports_inv,           --    reset_sink.reset_n
			islv_readdata    => eim_slave_to_avalon_master_0_avalon_master_readdata,    -- avalon_master.readdata
			islv_waitrequest => eim_slave_to_avalon_master_0_avalon_master_waitrequest, --              .waitrequest
			oslv_address     => eim_slave_to_avalon_master_0_avalon_master_address,     --              .address
			oslv_read        => eim_slave_to_avalon_master_0_avalon_master_read,        --              .read
			oslv_write       => eim_slave_to_avalon_master_0_avalon_master_write,       --              .write
			oslv_writedata   => eim_slave_to_avalon_master_0_avalon_master_writedata    --              .writedata
		);

	dacad5668_0 : component avalon_dacad5668_interface
		generic map (
			BASE_CLK           => 200000000,
			SCLK_FREQUENCY     => 10000000,
			INTERNAL_REFERENCE => '0',
			UNIQUE_ID          => "00010010011100000010000000000001"
		)
		port map (
			isl_clk             => altpll_0_c0_clk,                                                     --   clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                        --   reset_sink.reset_n
			osl_sclk            => dacad5668_0_conduit_end_osl_sclk,                                    --  conduit_end.export
			oslv_Ss             => dacad5668_0_conduit_end_oslv_Ss,                                     --             .export
			osl_mosi            => dacad5668_0_conduit_end_osl_mosi,                                    --             .export
			osl_LDAC_n          => dacad5668_0_conduit_end_osl_LDAC_n,                                  --             .export
			osl_CLR_n           => dacad5668_0_conduit_end_osl_CLR_n,                                   --             .export
			islv_avs_address    => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_address,     -- avalon_slave.address
			isl_avs_read        => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_read,        --             .read
			isl_avs_write       => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_write,       --             .write
			islv_avs_write_data => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_writedata,   --             .writedata
			oslv_avs_read_data  => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_readdata,    --             .readdata
			osl_avs_waitrequest => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest, --             .waitrequest
			islv_avs_byteenable => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_byteenable   --             .byteenable
		);

	fqd_interface_0 : component avalon_fqd_counter_interface
		generic map (
			number_of_fqds => 8,
			unique_id      => "00010010011100000110000000000001"
		)
		port map (
			oslv_avs_read_data  => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,    -- avalon_slave_0.readdata
			isl_avs_read        => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_read,        --               .read
			isl_avs_write       => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_write,       --               .write
			islv_avs_write_data => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,   --               .writedata
			islv_avs_address    => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_address,     --               .address
			osl_avs_waitrequest => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest, --               .waitrequest
			islv_avs_byteenable => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,  --               .byteenable
			isl_clk             => altpll_0_c0_clk,                                                           --     clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                              --     reset_sink.reset_n
			islv_enc_B          => fqd_interface_0_conduit_end_B,                                             --    conduit_end.export
			islv_enc_A          => fqd_interface_0_conduit_end_A                                              --               .export
		);

	gpio_block_0 : component cb20_gpio_block_0
		generic map (
			number_of_gpios => 9,
			unique_id       => "00010010011100000101000000000001"
		)
		port map (
			oslv_avs_read_data  => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,    -- avalon_slave_0.readdata
			islv_avs_address    => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address,     --               .address
			isl_avs_read        => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read,        --               .read
			isl_avs_write       => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write,       --               .write
			osl_avs_waitrequest => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest, --               .waitrequest
			islv_avs_write_data => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,   --               .writedata
			islv_avs_byteenable => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,  --               .byteenable
			isl_clk             => altpll_0_c0_clk,                                                        --     clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                           --     reset_sink.reset_n
			oslv_gpios          => gpio_block_0_conduit_end_export                                         --    conduit_end.export
		);

	pwm_interface_0 : component avalon_pwm_interface
		generic map (
			number_of_pwms => 4,
			base_clk       => 200000000,
			unique_id      => "00010010011100001100000000000001"
		)
		port map (
			oslv_avs_read_data  => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,    -- avalon_slave_0.readdata
			islv_avs_address    => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_address,     --               .address
			isl_avs_read        => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_read,        --               .read
			isl_avs_write       => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_write,       --               .write
			islv_avs_write_data => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,   --               .writedata
			osl_avs_waitrequest => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest, --               .waitrequest
			islv_avs_byteenable => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,  --               .byteenable
			isl_clk             => altpll_0_c0_clk,                                                           --     clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                              --     reset_sink.reset_n
			oslv_pwm            => pwm_interface_0_conduit_end_export                                         --    conduit_end.export
		);

	gpio_block_1 : component cb20_gpio_block_1
		generic map (
			number_of_gpios => 8,
			unique_id       => "00010010011100000101000000000010"
		)
		port map (
			oslv_avs_read_data  => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata,    -- avalon_slave_0.readdata
			islv_avs_address    => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_address,     --               .address
			isl_avs_read        => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_read,        --               .read
			isl_avs_write       => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_write,       --               .write
			osl_avs_waitrequest => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest, --               .waitrequest
			islv_avs_write_data => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata,   --               .writedata
			islv_avs_byteenable => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,  --               .byteenable
			isl_clk             => altpll_0_c0_clk,                                                        --     clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                           --     reset_sink.reset_n
			oslv_gpios          => gpio_block_1_conduit_end_export                                         --    conduit_end.export
		);

	watchdog_block_0 : component avalon_watchdog_interface
		generic map (
			base_clk  => 200000000,
			unique_id => "00010010011100010000000000000001"
		)
		port map (
			islv_avs_write_data => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,   -- avalon_slave_0.writedata
			oslv_avs_read_data  => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,    --               .readdata
			isl_avs_write       => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write,       --               .write
			isl_avs_read        => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read,        --               .read
			islv_avs_address    => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address,     --               .address
			osl_avs_waitrequest => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest, --               .waitrequest
			islv_avs_byteenable => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,  --               .byteenable
			isl_clk             => altpll_0_c0_clk,                                                            --     clock_sink.clk
			isl_reset_n         => rst_controller_001_reset_out_reset_ports_inv,                               --     reset_sink.reset_n
			osl_granted         => watchdog_block_0_wd_signals_granted,                                        --     wd_signals.export
			osl_watchdog_pwm    => watchdog_block_0_wd_signals_watchdog_pwm                                    --               .export
		);

	ppwa_block_0 : component avalon_ppwa_interface
		generic map (
			number_of_ppwas => 2,
			base_clk        => 200000000,
			unique_id       => "00010010011100001101000000000001"
		)
		port map (
			islv_avs_write_data     => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,   -- avalon_slave_0.writedata
			oslv_avs_read_data      => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,    --               .readdata
			islv_avs_address        => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address,     --               .address
			isl_avs_read            => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read,        --               .read
			isl_avs_write           => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write,       --               .write
			osl_avs_waitrequest     => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest, --               .waitrequest
			islv_avs_byteenable     => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,  --               .byteenable
			isl_clk                 => altpll_0_c0_clk,                                                        --     clock_sink.clk
			isl_reset_n             => rst_controller_001_reset_out_reset_ports_inv,                           --     reset_sink.reset_n
			islv_signals_to_measure => ppwa_block_0_conduit_end_export                                         --    conduit_end.export
		);

	eim_slave_to_avalon_master_0_avalon_master_translator : component altera_merlin_master_translator
		generic map (
			AV_ADDRESS_W                => 16,
			AV_DATA_W                   => 16,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 2,
			UAV_ADDRESS_W               => 17,
			UAV_BURSTCOUNT_W            => 2,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 2,
			AV_ADDRESS_SYMBOLS          => 0,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                               --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                            --                     reset.reset
			uav_address              => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => eim_slave_to_avalon_master_0_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => eim_slave_to_avalon_master_0_avalon_master_waitrequest,                                        --                          .waitrequest
			av_read                  => eim_slave_to_avalon_master_0_avalon_master_read,                                               --                          .read
			av_readdata              => eim_slave_to_avalon_master_0_avalon_master_readdata,                                           --                          .readdata
			av_write                 => eim_slave_to_avalon_master_0_avalon_master_write,                                              --                          .write
			av_writedata             => eim_slave_to_avalon_master_0_avalon_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                                           --               (terminated)
			av_byteenable            => "11",                                                                                          --               (terminated)
			av_beginbursttransfer    => '0',                                                                                           --               (terminated)
			av_begintransfer         => '0',                                                                                           --               (terminated)
			av_chipselect            => '0',                                                                                           --               (terminated)
			av_readdatavalid         => open,                                                                                          --               (terminated)
			av_lock                  => '0',                                                                                           --               (terminated)
			av_debugaccess           => '0',                                                                                           --               (terminated)
			uav_clken                => open,                                                                                          --               (terminated)
			av_clken                 => '1',                                                                                           --               (terminated)
			uav_response             => "00",                                                                                          --               (terminated)
			av_response              => open,                                                                                          --               (terminated)
			uav_writeresponserequest => open,                                                                                          --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                           --               (terminated)
			av_writeresponserequest  => '0',                                                                                           --               (terminated)
			av_writeresponsevalid    => open                                                                                           --               (terminated)
		);

	info_device_0_avalon_slave_translator : component cb20_info_device_0_avalon_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                       --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                    --                    reset.reset
			uav_address              => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => info_device_0_avalon_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => info_device_0_avalon_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => info_device_0_avalon_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => info_device_0_avalon_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => info_device_0_avalon_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => info_device_0_avalon_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => info_device_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                                  --              (terminated)
			av_burstcount            => open,                                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                                  --              (terminated)
			av_lock                  => open,                                                                                  --              (terminated)
			av_chipselect            => open,                                                                                  --              (terminated)
			av_clken                 => open,                                                                                  --              (terminated)
			uav_clken                => '0',                                                                                   --              (terminated)
			av_debugaccess           => open,                                                                                  --              (terminated)
			av_outputenable          => open,                                                                                  --              (terminated)
			uav_response             => open,                                                                                  --              (terminated)
			av_response              => "00",                                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                                    --              (terminated)
		);

	dacad5668_0_avalon_slave_translator : component cb20_info_device_0_avalon_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                     --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                  --                    reset.reset
			uav_address              => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => dacad5668_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                                --              (terminated)
			av_burstcount            => open,                                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                                --              (terminated)
			av_lock                  => open,                                                                                --              (terminated)
			av_chipselect            => open,                                                                                --              (terminated)
			av_clken                 => open,                                                                                --              (terminated)
			uav_clken                => '0',                                                                                 --              (terminated)
			av_debugaccess           => open,                                                                                --              (terminated)
			av_outputenable          => open,                                                                                --              (terminated)
			uav_response             => open,                                                                                --              (terminated)
			av_response              => "00",                                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                                  --              (terminated)
		);

	fqd_interface_0_avalon_slave_0_translator : component cb20_info_device_0_avalon_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                        --                    reset.reset
			uav_address              => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => fqd_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	gpio_block_0_avalon_slave_0_translator : component cb20_gpio_block_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                     --                    reset.reset
			uav_address              => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => gpio_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	pwm_interface_0_avalon_slave_0_translator : component cb20_pwm_interface_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 6,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                        --                    reset.reset
			uav_address              => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => pwm_interface_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	gpio_block_1_avalon_slave_0_translator : component cb20_gpio_block_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                     --                    reset.reset
			uav_address              => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => gpio_block_1_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	watchdog_block_0_avalon_slave_0_translator : component cb20_info_device_0_avalon_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                            --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                         --                    reset.reset
			uav_address              => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => watchdog_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                       --              (terminated)
			av_beginbursttransfer    => open,                                                                                       --              (terminated)
			av_burstcount            => open,                                                                                       --              (terminated)
			av_readdatavalid         => '0',                                                                                        --              (terminated)
			av_writebyteenable       => open,                                                                                       --              (terminated)
			av_lock                  => open,                                                                                       --              (terminated)
			av_chipselect            => open,                                                                                       --              (terminated)
			av_clken                 => open,                                                                                       --              (terminated)
			uav_clken                => '0',                                                                                        --              (terminated)
			av_debugaccess           => open,                                                                                       --              (terminated)
			av_outputenable          => open,                                                                                       --              (terminated)
			uav_response             => open,                                                                                       --              (terminated)
			av_response              => "00",                                                                                       --              (terminated)
			uav_writeresponserequest => '0',                                                                                        --              (terminated)
			uav_writeresponsevalid   => open,                                                                                       --              (terminated)
			av_writeresponserequest  => open,                                                                                       --              (terminated)
			av_writeresponsevalid    => '0'                                                                                         --              (terminated)
		);

	ppwa_block_0_avalon_slave_0_translator : component cb20_info_device_0_avalon_slave_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 17,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => altpll_0_c0_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                     --                    reset.reset
			uav_address              => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => ppwa_block_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 63,
			PKT_PROTECTION_L          => 61,
			PKT_BEGIN_BURST           => 52,
			PKT_BURSTWRAP_H           => 44,
			PKT_BURSTWRAP_L           => 44,
			PKT_BURST_SIZE_H          => 47,
			PKT_BURST_SIZE_L          => 45,
			PKT_BURST_TYPE_H          => 49,
			PKT_BURST_TYPE_L          => 48,
			PKT_BYTE_CNT_H            => 43,
			PKT_BYTE_CNT_L            => 41,
			PKT_ADDR_H                => 34,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 35,
			PKT_TRANS_POSTED          => 36,
			PKT_TRANS_WRITE           => 37,
			PKT_TRANS_READ            => 38,
			PKT_TRANS_LOCK            => 39,
			PKT_TRANS_EXCLUSIVE       => 40,
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_SRC_ID_H              => 56,
			PKT_SRC_ID_L              => 54,
			PKT_DEST_ID_H             => 59,
			PKT_DEST_ID_L             => 57,
			PKT_THREAD_ID_H           => 60,
			PKT_THREAD_ID_L           => 60,
			PKT_CACHE_H               => 67,
			PKT_CACHE_L               => 64,
			PKT_DATA_SIDEBAND_H       => 51,
			PKT_DATA_SIDEBAND_L       => 51,
			PKT_QOS_H                 => 53,
			PKT_QOS_L                 => 53,
			PKT_ADDR_SIDEBAND_H       => 50,
			PKT_ADDR_SIDEBAND_L       => 50,
			PKT_RESPONSE_STATUS_H     => 69,
			PKT_RESPONSE_STATUS_L     => 68,
			ST_DATA_W                 => 70,
			ST_CHANNEL_W              => 8,
			AV_BURSTCOUNT_W           => 2,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                        --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                     -- clk_reset.reset
			av_address              => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                                                 --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                                                  --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                                               --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                                         --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                                           --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                                                 --          .ready
			av_response             => open,                                                                                                   -- (terminated)
			av_writeresponserequest => '0',                                                                                                    -- (terminated)
			av_writeresponsevalid   => open                                                                                                    -- (terminated)
		);

	info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                 --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                              --       clk_reset.reset
			m0_address              => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_src_ready,                                                                         --              cp.ready
			cp_valid                => width_adapter_src_valid,                                                                         --                .valid
			cp_data                 => width_adapter_src_data,                                                                          --                .data
			cp_startofpacket        => width_adapter_src_startofpacket,                                                                 --                .startofpacket
			cp_endofpacket          => width_adapter_src_endofpacket,                                                                   --                .endofpacket
			cp_channel              => width_adapter_src_channel,                                                                       --                .channel
			rf_sink_ready           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                              --     (terminated)
		);

	info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                 --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                            -- (terminated)
			csr_read          => '0',                                                                                             -- (terminated)
			csr_write         => '0',                                                                                             -- (terminated)
			csr_readdata      => open,                                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                              -- (terminated)
			almost_full_data  => open,                                                                                            -- (terminated)
			almost_empty_data => open,                                                                                            -- (terminated)
			in_empty          => '0',                                                                                             -- (terminated)
			out_empty         => open,                                                                                            -- (terminated)
			in_error          => '0',                                                                                             -- (terminated)
			out_error         => open,                                                                                            -- (terminated)
			in_channel        => '0',                                                                                             -- (terminated)
			out_channel       => open                                                                                             -- (terminated)
		);

	dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                               --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_002_src_ready,                                                                   --              cp.ready
			cp_valid                => width_adapter_002_src_valid,                                                                   --                .valid
			cp_data                 => width_adapter_002_src_data,                                                                    --                .data
			cp_startofpacket        => width_adapter_002_src_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => width_adapter_002_src_endofpacket,                                                             --                .endofpacket
			cp_channel              => width_adapter_002_src_channel,                                                                 --                .channel
			rf_sink_ready           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                            --     (terminated)
		);

	dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                               --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                          -- (terminated)
			csr_read          => '0',                                                                                           -- (terminated)
			csr_write         => '0',                                                                                           -- (terminated)
			csr_readdata      => open,                                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                            -- (terminated)
			almost_full_data  => open,                                                                                          -- (terminated)
			almost_empty_data => open,                                                                                          -- (terminated)
			in_empty          => '0',                                                                                           -- (terminated)
			out_empty         => open,                                                                                          -- (terminated)
			in_error          => '0',                                                                                           -- (terminated)
			out_error         => open,                                                                                          -- (terminated)
			in_channel        => '0',                                                                                           -- (terminated)
			out_channel       => open                                                                                           -- (terminated)
		);

	fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                  --       clk_reset.reset
			m0_address              => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_004_src_ready,                                                                         --              cp.ready
			cp_valid                => width_adapter_004_src_valid,                                                                         --                .valid
			cp_data                 => width_adapter_004_src_data,                                                                          --                .data
			cp_startofpacket        => width_adapter_004_src_startofpacket,                                                                 --                .startofpacket
			cp_endofpacket          => width_adapter_004_src_endofpacket,                                                                   --                .endofpacket
			cp_channel              => width_adapter_004_src_channel,                                                                       --                .channel
			rf_sink_ready           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_006_src_ready,                                                                      --              cp.ready
			cp_valid                => width_adapter_006_src_valid,                                                                      --                .valid
			cp_data                 => width_adapter_006_src_data,                                                                       --                .data
			cp_startofpacket        => width_adapter_006_src_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => width_adapter_006_src_endofpacket,                                                                --                .endofpacket
			cp_channel              => width_adapter_006_src_channel,                                                                    --                .channel
			rf_sink_ready           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                  --       clk_reset.reset
			m0_address              => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_008_src_ready,                                                                         --              cp.ready
			cp_valid                => width_adapter_008_src_valid,                                                                         --                .valid
			cp_data                 => width_adapter_008_src_data,                                                                          --                .data
			cp_startofpacket        => width_adapter_008_src_startofpacket,                                                                 --                .startofpacket
			cp_endofpacket          => width_adapter_008_src_endofpacket,                                                                   --                .endofpacket
			cp_channel              => width_adapter_008_src_channel,                                                                       --                .channel
			rf_sink_ready           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_010_src_ready,                                                                      --              cp.ready
			cp_valid                => width_adapter_010_src_valid,                                                                      --                .valid
			cp_data                 => width_adapter_010_src_data,                                                                       --                .data
			cp_startofpacket        => width_adapter_010_src_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => width_adapter_010_src_endofpacket,                                                                --                .endofpacket
			cp_channel              => width_adapter_010_src_channel,                                                                    --                .channel
			rf_sink_ready           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                      --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_012_src_ready,                                                                          --              cp.ready
			cp_valid                => width_adapter_012_src_valid,                                                                          --                .valid
			cp_data                 => width_adapter_012_src_data,                                                                           --                .data
			cp_startofpacket        => width_adapter_012_src_startofpacket,                                                                  --                .startofpacket
			cp_endofpacket          => width_adapter_012_src_endofpacket,                                                                    --                .endofpacket
			cp_channel              => width_adapter_012_src_channel,                                                                        --                .channel
			rf_sink_ready           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                 --     (terminated)
			m0_writeresponserequest => open,                                                                                                 --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                   --     (terminated)
		);

	watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                      --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                 -- (terminated)
			csr_read          => '0',                                                                                                  -- (terminated)
			csr_write         => '0',                                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                   -- (terminated)
			almost_full_data  => open,                                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                                 -- (terminated)
			in_empty          => '0',                                                                                                  -- (terminated)
			out_empty         => open,                                                                                                 -- (terminated)
			in_error          => '0',                                                                                                  -- (terminated)
			out_error         => open,                                                                                                 -- (terminated)
			in_channel        => '0',                                                                                                  -- (terminated)
			out_channel       => open                                                                                                  -- (terminated)
		);

	ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 52,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 53,
			PKT_TRANS_POSTED          => 54,
			PKT_TRANS_WRITE           => 55,
			PKT_TRANS_READ            => 56,
			PKT_TRANS_LOCK            => 57,
			PKT_SRC_ID_H              => 74,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 77,
			PKT_DEST_ID_L             => 75,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 62,
			PKT_BYTE_CNT_H            => 61,
			PKT_BYTE_CNT_L            => 59,
			PKT_PROTECTION_H          => 81,
			PKT_PROTECTION_L          => 79,
			PKT_RESPONSE_STATUS_H     => 87,
			PKT_RESPONSE_STATUS_L     => 86,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 88,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => altpll_0_c0_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_014_src_ready,                                                                      --              cp.ready
			cp_valid                => width_adapter_014_src_valid,                                                                      --                .valid
			cp_data                 => width_adapter_014_src_data,                                                                       --                .data
			cp_startofpacket        => width_adapter_014_src_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => width_adapter_014_src_endofpacket,                                                                --                .endofpacket
			cp_channel              => width_adapter_014_src_channel,                                                                    --                .channel
			rf_sink_ready           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 89,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => altpll_0_c0_clk,                                                                                  --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	addr_router : component cb20_addr_router
		port map (
			sink_ready         => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => eim_slave_to_avalon_master_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                                  --       src.ready
			src_valid          => addr_router_src_valid,                                                                                  --          .valid
			src_data           => addr_router_src_data,                                                                                   --          .data
			src_channel        => addr_router_src_channel,                                                                                --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                                          --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                             --          .endofpacket
		);

	id_router : component cb20_id_router
		port map (
			sink_ready         => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => info_device_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                   --       src.ready
			src_valid          => id_router_src_valid,                                                                   --          .valid
			src_data           => id_router_src_data,                                                                    --          .data
			src_channel        => id_router_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                              --          .endofpacket
		);

	id_router_001 : component cb20_id_router
		port map (
			sink_ready         => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => dacad5668_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                             --       src.ready
			src_valid          => id_router_001_src_valid,                                                             --          .valid
			src_data           => id_router_001_src_data,                                                              --          .data
			src_channel        => id_router_001_src_channel,                                                           --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                        --          .endofpacket
		);

	id_router_002 : component cb20_id_router
		port map (
			sink_ready         => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => fqd_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                   --       src.ready
			src_valid          => id_router_002_src_valid,                                                                   --          .valid
			src_data           => id_router_002_src_data,                                                                    --          .data
			src_channel        => id_router_002_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                              --          .endofpacket
		);

	id_router_003 : component cb20_id_router
		port map (
			sink_ready         => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => gpio_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                                --       src.ready
			src_valid          => id_router_003_src_valid,                                                                --          .valid
			src_data           => id_router_003_src_data,                                                                 --          .data
			src_channel        => id_router_003_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                           --          .endofpacket
		);

	id_router_004 : component cb20_id_router
		port map (
			sink_ready         => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pwm_interface_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                   --       src.ready
			src_valid          => id_router_004_src_valid,                                                                   --          .valid
			src_data           => id_router_004_src_data,                                                                    --          .data
			src_channel        => id_router_004_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                              --          .endofpacket
		);

	id_router_005 : component cb20_id_router
		port map (
			sink_ready         => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => gpio_block_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                                --       src.ready
			src_valid          => id_router_005_src_valid,                                                                --          .valid
			src_data           => id_router_005_src_data,                                                                 --          .data
			src_channel        => id_router_005_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                           --          .endofpacket
		);

	id_router_006 : component cb20_id_router
		port map (
			sink_ready         => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => watchdog_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                    --       src.ready
			src_valid          => id_router_006_src_valid,                                                                    --          .valid
			src_data           => id_router_006_src_data,                                                                     --          .data
			src_channel        => id_router_006_src_channel,                                                                  --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                            --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                               --          .endofpacket
		);

	id_router_007 : component cb20_id_router
		port map (
			sink_ready         => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ppwa_block_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => altpll_0_c0_clk,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                                --       src.ready
			src_valid          => id_router_007_src_valid,                                                                --          .valid
			src_data           => id_router_007_src_data,                                                                 --          .data
			src_channel        => id_router_007_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                           --          .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => altpll_0_c0_clk,                    --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component cb20_cmd_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                    --       clk.clk
			reset              => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sink_ready         => addr_router_src_ready,              --      sink.ready
			sink_channel       => addr_router_src_channel,            --          .channel
			sink_data          => addr_router_src_data,               --          .data
			sink_startofpacket => addr_router_src_startofpacket,      --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,        --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,              --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,          --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,          --          .valid
			src0_data          => cmd_xbar_demux_src0_data,           --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,        --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket,  --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,    --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,          --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,          --          .valid
			src1_data          => cmd_xbar_demux_src1_data,           --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,        --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket,  --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,    --          .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,          --      src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,          --          .valid
			src2_data          => cmd_xbar_demux_src2_data,           --          .data
			src2_channel       => cmd_xbar_demux_src2_channel,        --          .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket,  --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket,    --          .endofpacket
			src3_ready         => cmd_xbar_demux_src3_ready,          --      src3.ready
			src3_valid         => cmd_xbar_demux_src3_valid,          --          .valid
			src3_data          => cmd_xbar_demux_src3_data,           --          .data
			src3_channel       => cmd_xbar_demux_src3_channel,        --          .channel
			src3_startofpacket => cmd_xbar_demux_src3_startofpacket,  --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_src3_endofpacket,    --          .endofpacket
			src4_ready         => cmd_xbar_demux_src4_ready,          --      src4.ready
			src4_valid         => cmd_xbar_demux_src4_valid,          --          .valid
			src4_data          => cmd_xbar_demux_src4_data,           --          .data
			src4_channel       => cmd_xbar_demux_src4_channel,        --          .channel
			src4_startofpacket => cmd_xbar_demux_src4_startofpacket,  --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_src4_endofpacket,    --          .endofpacket
			src5_ready         => cmd_xbar_demux_src5_ready,          --      src5.ready
			src5_valid         => cmd_xbar_demux_src5_valid,          --          .valid
			src5_data          => cmd_xbar_demux_src5_data,           --          .data
			src5_channel       => cmd_xbar_demux_src5_channel,        --          .channel
			src5_startofpacket => cmd_xbar_demux_src5_startofpacket,  --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_src5_endofpacket,    --          .endofpacket
			src6_ready         => cmd_xbar_demux_src6_ready,          --      src6.ready
			src6_valid         => cmd_xbar_demux_src6_valid,          --          .valid
			src6_data          => cmd_xbar_demux_src6_data,           --          .data
			src6_channel       => cmd_xbar_demux_src6_channel,        --          .channel
			src6_startofpacket => cmd_xbar_demux_src6_startofpacket,  --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_src6_endofpacket,    --          .endofpacket
			src7_ready         => cmd_xbar_demux_src7_ready,          --      src7.ready
			src7_valid         => cmd_xbar_demux_src7_valid,          --          .valid
			src7_data          => cmd_xbar_demux_src7_data,           --          .data
			src7_channel       => cmd_xbar_demux_src7_channel,        --          .channel
			src7_startofpacket => cmd_xbar_demux_src7_startofpacket,  --          .startofpacket
			src7_endofpacket   => cmd_xbar_demux_src7_endofpacket     --          .endofpacket
		);

	rsp_xbar_demux : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,         --      sink.ready
			sink_channel       => width_adapter_001_src_channel,       --          .channel
			sink_data          => width_adapter_001_src_data,          --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket, --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,   --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,         --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,           --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,           --          .valid
			src0_data          => rsp_xbar_demux_src0_data,            --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,         --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket,   --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket      --          .endofpacket
		);

	rsp_xbar_demux_001 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_003_src_ready,           --      sink.ready
			sink_channel       => width_adapter_003_src_channel,         --          .channel
			sink_data          => width_adapter_003_src_data,            --          .data
			sink_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_003_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_005_src_ready,           --      sink.ready
			sink_channel       => width_adapter_005_src_channel,         --          .channel
			sink_data          => width_adapter_005_src_data,            --          .data
			sink_startofpacket => width_adapter_005_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_005_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_005_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_007_src_ready,           --      sink.ready
			sink_channel       => width_adapter_007_src_channel,         --          .channel
			sink_data          => width_adapter_007_src_data,            --          .data
			sink_startofpacket => width_adapter_007_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_007_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_007_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_009_src_ready,           --      sink.ready
			sink_channel       => width_adapter_009_src_channel,         --          .channel
			sink_data          => width_adapter_009_src_data,            --          .data
			sink_startofpacket => width_adapter_009_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_009_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_009_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_011_src_ready,           --      sink.ready
			sink_channel       => width_adapter_011_src_channel,         --          .channel
			sink_data          => width_adapter_011_src_data,            --          .data
			sink_startofpacket => width_adapter_011_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_011_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_011_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_013_src_ready,           --      sink.ready
			sink_channel       => width_adapter_013_src_channel,         --          .channel
			sink_data          => width_adapter_013_src_data,            --          .data
			sink_startofpacket => width_adapter_013_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_013_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_013_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component cb20_rsp_xbar_demux
		port map (
			clk                => altpll_0_c0_clk,                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_015_src_ready,           --      sink.ready
			sink_channel       => width_adapter_015_src_channel,         --          .channel
			sink_data          => width_adapter_015_src_data,            --          .data
			sink_startofpacket => width_adapter_015_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_015_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_015_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component cb20_rsp_xbar_mux
		port map (
			clk                 => altpll_0_c0_clk,                       --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready         => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data          => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                    --       clk.clk
			reset                => rst_controller_001_reset_out_reset, -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src0_valid,          --      sink.valid
			in_channel           => cmd_xbar_demux_src0_channel,        --          .channel
			in_startofpacket     => cmd_xbar_demux_src0_startofpacket,  --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src0_endofpacket,    --          .endofpacket
			in_ready             => cmd_xbar_demux_src0_ready,          --          .ready
			in_data              => cmd_xbar_demux_src0_data,           --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_src_valid,                 --      sink.valid
			in_channel           => id_router_src_channel,               --          .channel
			in_startofpacket     => id_router_src_startofpacket,         --          .startofpacket
			in_endofpacket       => id_router_src_endofpacket,           --          .endofpacket
			in_ready             => id_router_src_ready,                 --          .ready
			in_data              => id_router_src_data,                  --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_002 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src1_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src1_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src1_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src1_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src1_ready,           --          .ready
			in_data              => cmd_xbar_demux_src1_data,            --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_002_src_data,          --          .data
			out_channel          => width_adapter_002_src_channel,       --          .channel
			out_valid            => width_adapter_002_src_valid,         --          .valid
			out_ready            => width_adapter_002_src_ready,         --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_003 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_001_src_valid,             --      sink.valid
			in_channel           => id_router_001_src_channel,           --          .channel
			in_startofpacket     => id_router_001_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_001_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_001_src_ready,             --          .ready
			in_data              => id_router_001_src_data,              --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_003_src_data,          --          .data
			out_channel          => width_adapter_003_src_channel,       --          .channel
			out_valid            => width_adapter_003_src_valid,         --          .valid
			out_ready            => width_adapter_003_src_ready,         --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_004 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src2_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src2_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src2_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src2_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src2_ready,           --          .ready
			in_data              => cmd_xbar_demux_src2_data,            --          .data
			out_endofpacket      => width_adapter_004_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_004_src_data,          --          .data
			out_channel          => width_adapter_004_src_channel,       --          .channel
			out_valid            => width_adapter_004_src_valid,         --          .valid
			out_ready            => width_adapter_004_src_ready,         --          .ready
			out_startofpacket    => width_adapter_004_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_005 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_002_src_valid,             --      sink.valid
			in_channel           => id_router_002_src_channel,           --          .channel
			in_startofpacket     => id_router_002_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_002_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_002_src_ready,             --          .ready
			in_data              => id_router_002_src_data,              --          .data
			out_endofpacket      => width_adapter_005_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_005_src_data,          --          .data
			out_channel          => width_adapter_005_src_channel,       --          .channel
			out_valid            => width_adapter_005_src_valid,         --          .valid
			out_ready            => width_adapter_005_src_ready,         --          .ready
			out_startofpacket    => width_adapter_005_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_006 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src3_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src3_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src3_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src3_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src3_ready,           --          .ready
			in_data              => cmd_xbar_demux_src3_data,            --          .data
			out_endofpacket      => width_adapter_006_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_006_src_data,          --          .data
			out_channel          => width_adapter_006_src_channel,       --          .channel
			out_valid            => width_adapter_006_src_valid,         --          .valid
			out_ready            => width_adapter_006_src_ready,         --          .ready
			out_startofpacket    => width_adapter_006_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_007 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_003_src_valid,             --      sink.valid
			in_channel           => id_router_003_src_channel,           --          .channel
			in_startofpacket     => id_router_003_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_003_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_003_src_ready,             --          .ready
			in_data              => id_router_003_src_data,              --          .data
			out_endofpacket      => width_adapter_007_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_007_src_data,          --          .data
			out_channel          => width_adapter_007_src_channel,       --          .channel
			out_valid            => width_adapter_007_src_valid,         --          .valid
			out_ready            => width_adapter_007_src_ready,         --          .ready
			out_startofpacket    => width_adapter_007_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_008 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src4_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src4_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src4_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src4_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src4_ready,           --          .ready
			in_data              => cmd_xbar_demux_src4_data,            --          .data
			out_endofpacket      => width_adapter_008_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_008_src_data,          --          .data
			out_channel          => width_adapter_008_src_channel,       --          .channel
			out_valid            => width_adapter_008_src_valid,         --          .valid
			out_ready            => width_adapter_008_src_ready,         --          .ready
			out_startofpacket    => width_adapter_008_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_009 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_004_src_valid,             --      sink.valid
			in_channel           => id_router_004_src_channel,           --          .channel
			in_startofpacket     => id_router_004_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_004_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_004_src_ready,             --          .ready
			in_data              => id_router_004_src_data,              --          .data
			out_endofpacket      => width_adapter_009_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_009_src_data,          --          .data
			out_channel          => width_adapter_009_src_channel,       --          .channel
			out_valid            => width_adapter_009_src_valid,         --          .valid
			out_ready            => width_adapter_009_src_ready,         --          .ready
			out_startofpacket    => width_adapter_009_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_010 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src5_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src5_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src5_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src5_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src5_ready,           --          .ready
			in_data              => cmd_xbar_demux_src5_data,            --          .data
			out_endofpacket      => width_adapter_010_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_010_src_data,          --          .data
			out_channel          => width_adapter_010_src_channel,       --          .channel
			out_valid            => width_adapter_010_src_valid,         --          .valid
			out_ready            => width_adapter_010_src_ready,         --          .ready
			out_startofpacket    => width_adapter_010_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_011 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_005_src_valid,             --      sink.valid
			in_channel           => id_router_005_src_channel,           --          .channel
			in_startofpacket     => id_router_005_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_005_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_005_src_ready,             --          .ready
			in_data              => id_router_005_src_data,              --          .data
			out_endofpacket      => width_adapter_011_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_011_src_data,          --          .data
			out_channel          => width_adapter_011_src_channel,       --          .channel
			out_valid            => width_adapter_011_src_valid,         --          .valid
			out_ready            => width_adapter_011_src_ready,         --          .ready
			out_startofpacket    => width_adapter_011_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_012 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src6_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src6_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src6_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src6_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src6_ready,           --          .ready
			in_data              => cmd_xbar_demux_src6_data,            --          .data
			out_endofpacket      => width_adapter_012_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_012_src_data,          --          .data
			out_channel          => width_adapter_012_src_channel,       --          .channel
			out_valid            => width_adapter_012_src_valid,         --          .valid
			out_ready            => width_adapter_012_src_ready,         --          .ready
			out_startofpacket    => width_adapter_012_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_013 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_006_src_valid,             --      sink.valid
			in_channel           => id_router_006_src_channel,           --          .channel
			in_startofpacket     => id_router_006_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_006_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_006_src_ready,             --          .ready
			in_data              => id_router_006_src_data,              --          .data
			out_endofpacket      => width_adapter_013_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_013_src_data,          --          .data
			out_channel          => width_adapter_013_src_channel,       --          .channel
			out_valid            => width_adapter_013_src_valid,         --          .valid
			out_ready            => width_adapter_013_src_ready,         --          .ready
			out_startofpacket    => width_adapter_013_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_014 : component cb20_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 34,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 43,
			IN_PKT_BYTE_CNT_L             => 41,
			IN_PKT_TRANS_COMPRESSED_READ  => 35,
			IN_PKT_BURSTWRAP_H            => 44,
			IN_PKT_BURSTWRAP_L            => 44,
			IN_PKT_BURST_SIZE_H           => 47,
			IN_PKT_BURST_SIZE_L           => 45,
			IN_PKT_RESPONSE_STATUS_H      => 69,
			IN_PKT_RESPONSE_STATUS_L      => 68,
			IN_PKT_TRANS_EXCLUSIVE        => 40,
			IN_PKT_BURST_TYPE_H           => 49,
			IN_PKT_BURST_TYPE_L           => 48,
			IN_ST_DATA_W                  => 70,
			OUT_PKT_ADDR_H                => 52,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 61,
			OUT_PKT_BYTE_CNT_L            => 59,
			OUT_PKT_TRANS_COMPRESSED_READ => 53,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 87,
			OUT_PKT_RESPONSE_STATUS_L     => 86,
			OUT_PKT_TRANS_EXCLUSIVE       => 58,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 88,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src7_valid,           --      sink.valid
			in_channel           => cmd_xbar_demux_src7_channel,         --          .channel
			in_startofpacket     => cmd_xbar_demux_src7_startofpacket,   --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src7_endofpacket,     --          .endofpacket
			in_ready             => cmd_xbar_demux_src7_ready,           --          .ready
			in_data              => cmd_xbar_demux_src7_data,            --          .data
			out_endofpacket      => width_adapter_014_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_014_src_data,          --          .data
			out_channel          => width_adapter_014_src_channel,       --          .channel
			out_valid            => width_adapter_014_src_valid,         --          .valid
			out_ready            => width_adapter_014_src_ready,         --          .ready
			out_startofpacket    => width_adapter_014_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_015 : component cb20_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 52,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 61,
			IN_PKT_BYTE_CNT_L             => 59,
			IN_PKT_TRANS_COMPRESSED_READ  => 53,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 62,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 87,
			IN_PKT_RESPONSE_STATUS_L      => 86,
			IN_PKT_TRANS_EXCLUSIVE        => 58,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 88,
			OUT_PKT_ADDR_H                => 34,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 43,
			OUT_PKT_BYTE_CNT_L            => 41,
			OUT_PKT_TRANS_COMPRESSED_READ => 35,
			OUT_PKT_BURST_SIZE_H          => 47,
			OUT_PKT_BURST_SIZE_L          => 45,
			OUT_PKT_RESPONSE_STATUS_H     => 69,
			OUT_PKT_RESPONSE_STATUS_L     => 68,
			OUT_PKT_TRANS_EXCLUSIVE       => 40,
			OUT_PKT_BURST_TYPE_H          => 49,
			OUT_PKT_BURST_TYPE_L          => 48,
			OUT_ST_DATA_W                 => 70,
			ST_CHANNEL_W                  => 8,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => altpll_0_c0_clk,                     --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_007_src_valid,             --      sink.valid
			in_channel           => id_router_007_src_channel,           --          .channel
			in_startofpacket     => id_router_007_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_007_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_007_src_ready,             --          .ready
			in_data              => id_router_007_src_data,              --          .data
			out_endofpacket      => width_adapter_015_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_015_src_data,          --          .data
			out_channel          => width_adapter_015_src_channel,       --          .channel
			out_valid            => width_adapter_015_src_valid,         --          .valid
			out_ready            => width_adapter_015_src_ready,         --          .ready
			out_startofpacket    => width_adapter_015_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of cb20
